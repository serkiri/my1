library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity my1_top is
	port(
		CLK_20			: in std_logic;
		CLK_20_ALT		: in std_logic
	);
  
end my1_top;

architecture rtl of my1_top is

begin

end rtl;
